module draw_screen (x, y, objects, char_x, char_y, rgb, state);
	parameter object_num = 5;
	parameter char_width = 11;
	parameter char_height = 18;
	input logic [9:0] x;
	input logic [8:0] y;
	input logic [43:0] objects [object_num-1:0];
	input logic [9:0] char_x;
	input logic [8:0] char_y;
	output logic [23:0] rgb;
	input logic state;
	integer i;
	
	logic in_char;
	
	assign in_char = (x>=char_x)&(y>=char_y)&(x<=(char_x+char_width))&(y<=(char_y+char_height));
	always_comb begin
		rgb=0;
		for (i=0; i<object_num; i++) begin
			if ((objects[i][43:33]<=x)&(objects[i][32:22]<=y)&(objects[i][21:11]>=x)&(objects[i][10:0]>=y)) begin
				rgb = '1;
			end
		end
		if (in_char) begin
			case(state)
				1'b1: rgb = character[(y-char_y)/2][(x-char_x)/2];
				1'b0: rgb = character_jump[(y-char_y)/2][(x-char_x)/2];
			endcase
		end
	end //always_comb
	logic [23:0] character [char_height/2-1:0][char_width/2-1:0];
	always_comb begin
		character[0][0] = 24'b000000000000000000000000;
		character[0][1] = 24'b000000000000000000000000;
		character[0][2] = 24'b000000000000000000000000;
		character[0][3] = 24'b000000000000000000000000;
		character[0][4] = 24'b111111111111111111111111;
		character[0][5] = 24'b111111111111111111111111;
		character[0][6] = 24'b111111111111111111111111;
		character[0][7] = 24'b000000000000000000000000;
		character[0][8] = 24'b000000000000000000000000;
		character[0][9] = 24'b000000000000000000000000;
		character[0][10] = 24'b000000000000000000000000;
		character[1][0] = 24'b000000000000000000000000;
		character[1][1] = 24'b000000000000000000000000;
		character[1][2] = 24'b000000000000000000000000;
		character[1][3] = 24'b111111111111111111111111;
		character[1][4] = 24'b111111111010001110110001;
		character[1][5] = 24'b111111111010001110110001;
		character[1][6] = 24'b111111111010001110110001;
		character[1][7] = 24'b111111111111111111111111;
		character[1][8] = 24'b000000000000000000000000;
		character[1][9] = 24'b000000000000000000000000;
		character[1][10] = 24'b000000000000000000000000;
		character[2][0] = 24'b000000000000000000000000;
		character[2][1] = 24'b000000000000000000000000;
		character[2][2] = 24'b000000000000000000000000;
		character[2][3] = 24'b111111111010001110110001;
		character[2][4] = 24'b111111111010001110110001;
		character[2][5] = 24'b111111111010001110110001;
		character[2][6] = 24'b111111111010001110110001;
		character[2][7] = 24'b111111111010001110110001;
		character[2][8] = 24'b000000000000000000000000;
		character[2][9] = 24'b000000000000000000000000;
		character[2][10] = 24'b000000000000000000000000;
		character[3][0] = 24'b000000000000000000000000;
		character[3][1] = 24'b000000000000000000000000;
		character[3][2] = 24'b000000000000000000000000;
		character[3][3] = 24'b111111111010001110110001;
		character[3][4] = 24'b000000000000000000000000;
		character[3][5] = 24'b111111111010001110110001;
		character[3][6] = 24'b000000000000000000000000;
		character[3][7] = 24'b111111111010001110110001;
		character[3][8] = 24'b000000000000000000000000;
		character[3][9] = 24'b000000000000000000000000;
		character[3][10] = 24'b000000000000000000000000;
		character[4][0] = 24'b000000000000000000000000;
		character[4][1] = 24'b000000000000000000000000;
		character[4][2] = 24'b000000000000000000000000;
		character[4][3] = 24'b111111111010001110110001;
		character[4][4] = 24'b111111111010001110110001;
		character[4][5] = 24'b111111111010001110110001;
		character[4][6] = 24'b111111111010001110110001;
		character[4][7] = 24'b111111111010001110110001;
		character[4][8] = 24'b000000000000000000000000;
		character[4][9] = 24'b000000000000000000000000;
		character[4][10] = 24'b000000000000000000000000;
		character[5][0] = 24'b000000000000000000000000;
		character[5][1] = 24'b000000000000000000000000;
		character[5][2] = 24'b000000000000000000000000;
		character[5][3] = 24'b111111111010001110110001;
		character[5][4] = 24'b111111111010001110110001;
		character[5][5] = 24'b111111111010001110110001;
		character[5][6] = 24'b111111111010001110110001;
		character[5][7] = 24'b111111111010001110110001;
		character[5][8] = 24'b000000000000000000000000;
		character[5][9] = 24'b000000000000000000000000;
		character[5][10] = 24'b000000000000000000000000;
		character[6][0] = 24'b000000000000000000000000;
		character[6][1] = 24'b000000000000000000000000;
		character[6][2] = 24'b000000000000000000000000;
		character[6][3] = 24'b000000000000000000000000;
		character[6][4] = 24'b111111111010001110110001;
		character[6][5] = 24'b111111111010001110110001;
		character[6][6] = 24'b111111111010001110110001;
		character[6][7] = 24'b000000000000000000000000;
		character[6][8] = 24'b000000000000000000000000;
		character[6][9] = 24'b000000000000000000000000;
		character[6][10] = 24'b000000000000000000000000;
		character[7][0] = 24'b000000000000000000000000;
		character[7][1] = 24'b111111111010001110110001;
		character[7][2] = 24'b111111111111111111111111;
		character[7][3] = 24'b111111111010001110110001;
		character[7][4] = 24'b111111111010001110110001;
		character[7][5] = 24'b111111111010001110110001;
		character[7][6] = 24'b111111111010001110110001;
		character[7][7] = 24'b111111111010001110110001;
		character[7][8] = 24'b111111111111111111111111;
		character[7][9] = 24'b111111111010001110110001;
		character[7][10] = 24'b000000000000000000000000;
		character[8][0] = 24'b111111111010001110110001;
		character[8][1] = 24'b111111111010001110110001;
		character[8][2] = 24'b111111111111111111111111;
		character[8][3] = 24'b111111111111111111111111;
		character[8][4] = 24'b111111111010001110110001;
		character[8][5] = 24'b111111111010001110110001;
		character[8][6] = 24'b111111111010001110110001;
		character[8][7] = 24'b111111111111111111111111;
		character[8][8] = 24'b111111111111111111111111;
		character[8][9] = 24'b111111111010001110110001;
		character[8][10] = 24'b111111111010001110110001;
		character[9][0] = 24'b111111111010001110110001;
		character[9][1] = 24'b111111111010001110110001;
		character[9][2] = 24'b111111111111111111111111;
		character[9][3] = 24'b111111111111111111111111;
		character[9][4] = 24'b111111111111111111111111;
		character[9][5] = 24'b111111111010001110110001;
		character[9][6] = 24'b111111111111111111111111;
		character[9][7] = 24'b111111111111111111111111;
		character[9][8] = 24'b111111111111111111111111;
		character[9][9] = 24'b111111111010001110110001;
		character[9][10] = 24'b111111111010001110110001;
		character[10][0] = 24'b111111111010001110110001;
		character[10][1] = 24'b111111111010001110110001;
		character[10][2] = 24'b000000000000000000000000;
		character[10][3] = 24'b111111111111111111111111;
		character[10][4] = 24'b111111111111111111111111;
		character[10][5] = 24'b111111111111111111111111;
		character[10][6] = 24'b111111111111111111111111;
		character[10][7] = 24'b111111111111111111111111;
		character[10][8] = 24'b000000000000000000000000;
		character[10][9] = 24'b111111111010001110110001;
		character[10][10] = 24'b111111111010001110110001;
		character[11][0] = 24'b111111111010001110110001;
		character[11][1] = 24'b111111111010001110110001;
		character[11][2] = 24'b000000000000000000000000;
		character[11][3] = 24'b111111111111111111111111;
		character[11][4] = 24'b111111111111111111111111;
		character[11][5] = 24'b111111111111111111111111;
		character[11][6] = 24'b111111111111111111111111;
		character[11][7] = 24'b111111111111111111111111;
		character[11][8] = 24'b000000000000000000000000;
		character[11][9] = 24'b111111111010001110110001;
		character[11][10] = 24'b111111111010001110110001;
		character[12][0] = 24'b111111111010001110110001;
		character[12][1] = 24'b111111111010001110110001;
		character[12][2] = 24'b000000000000000000000000;
		character[12][3] = 24'b111111111111111111111111;
		character[12][4] = 24'b111111111111111111111111;
		character[12][5] = 24'b111111111111111111111111;
		character[12][6] = 24'b111111111111111111111111;
		character[12][7] = 24'b111111111111111111111111;
		character[12][8] = 24'b000000000000000000000000;
		character[12][9] = 24'b111111111010001110110001;
		character[12][10] = 24'b111111111010001110110001;
		character[13][0] = 24'b111111111111001000000000;
		character[13][1] = 24'b111111111010001110110001;
		character[13][2] = 24'b000000000000000000000000;
		character[13][3] = 24'b111111111111111111111111;
		character[13][4] = 24'b111111111111111111111111;
		character[13][5] = 24'b111111111111111111111111;
		character[13][6] = 24'b111111111111111111111111;
		character[13][7] = 24'b111111111111111111111111;
		character[13][8] = 24'b000000000000000000000000;
		character[13][9] = 24'b111111111010001110110001;
		character[13][10] = 24'b111111111111001000000000;
		character[14][0] = 24'b000000000000000000000000;
		character[14][1] = 24'b000000000000000000000000;
		character[14][2] = 24'b000000000000000000000000;
		character[14][3] = 24'b111111111111111111111111;
		character[14][4] = 24'b111111111111111111111111;
		character[14][5] = 24'b111111111111111111111111;
		character[14][6] = 24'b111111111111111111111111;
		character[14][7] = 24'b111111111111111111111111;
		character[14][8] = 24'b000000000000000000000000;
		character[14][9] = 24'b000000000000000000000000;
		character[14][10] = 24'b000000000000000000000000;
		character[15][0] = 24'b000000000000000000000000;
		character[15][1] = 24'b000000000000000000000000;
		character[15][2] = 24'b000000000000000000000000;
		character[15][3] = 24'b111111111111111111111111;
		character[15][4] = 24'b111111111111111111111111;
		character[15][5] = 24'b000000000000000000000000;
		character[15][6] = 24'b111111111111111111111111;
		character[15][7] = 24'b111111111111111111111111;
		character[15][8] = 24'b000000000000000000000000;
		character[15][9] = 24'b000000000000000000000000;
		character[15][10] = 24'b000000000000000000000000;
		character[16][0] = 24'b000000000000000000000000;
		character[16][1] = 24'b000000000000000000000000;
		character[16][2] = 24'b111111110111111000000000;
		character[16][3] = 24'b111111110111111000000000;
		character[16][4] = 24'b111111110111111000000000;
		character[16][5] = 24'b000000000000000000000000;
		character[16][6] = 24'b111111110111111000000000;
		character[16][7] = 24'b111111110111111000000000;
		character[16][8] = 24'b111111110111111000000000;
		character[16][9] = 24'b000000000000000000000000;
		character[16][10] = 24'b000000000000000000000000;
		character[17][0] = 24'b000000000000000000000000;
		character[17][1] = 24'b000000000000000000000000;
		character[17][2] = 24'b111111110111111000000000;
		character[17][3] = 24'b111111110111111000000000;
		character[17][4] = 24'b111111110111111000000000;
		character[17][5] = 24'b000000000000000000000000;
		character[17][6] = 24'b111111110111111000000000;
		character[17][7] = 24'b111111110111111000000000;
		character[17][8] = 24'b111111110111111000000000;
		character[17][9] = 24'b000000000000000000000000;
		character[17][10] = 24'b000000000000000000000000;
	end
	
	logic [23:0] character_jump [char_height/2-1:0][char_width/2-1:0];
	always_comb begin
		character_jump[0][0] = 24'b000000000000000000000000;
		character_jump[0][1] = 24'b000000000000000000000000;
		character_jump[0][2] = 24'b000000000000000000000000;
		character_jump[0][3] = 24'b000000000000000000000000;
		character_jump[0][4] = 24'b111111111111111111111111;
		character_jump[0][5] = 24'b111111111111111111111111;
		character_jump[0][6] = 24'b111111111111111111111111;
		character_jump[0][7] = 24'b000000000000000000000000;
		character_jump[0][8] = 24'b000000000000000000000000;
		character_jump[0][9] = 24'b000000000000000000000000;
		character_jump[0][10] = 24'b000000000000000000000000;
		character_jump[1][0] = 24'b000000000000000000000000;
		character_jump[1][1] = 24'b000000000000000000000000;
		character_jump[1][2] = 24'b000000000000000000000000;
		character_jump[1][3] = 24'b111111111111111111111111;
		character_jump[1][4] = 24'b111111111010001110110001;
		character_jump[1][5] = 24'b111111111010001110110001;
		character_jump[1][6] = 24'b111111111010001110110001;
		character_jump[1][7] = 24'b111111111111111111111111;
		character_jump[1][8] = 24'b000000000000000000000000;
		character_jump[1][9] = 24'b000000000000000000000000;
		character_jump[1][10] = 24'b000000000000000000000000;
		character_jump[2][0] = 24'b000000000000000000000000;
		character_jump[2][1] = 24'b000000000000000000000000;
		character_jump[2][2] = 24'b000000000000000000000000;
		character_jump[2][3] = 24'b111111111010001110110001;
		character_jump[2][4] = 24'b111111111010001110110001;
		character_jump[2][5] = 24'b111111111010001110110001;
		character_jump[2][6] = 24'b111111111010001110110001;
		character_jump[2][7] = 24'b111111111010001110110001;
		character_jump[2][8] = 24'b000000000000000000000000;
		character_jump[2][9] = 24'b000000000000000000000000;
		character_jump[2][10] = 24'b000000000000000000000000;
		character_jump[3][0] = 24'b111111111111001000000000;
		character_jump[3][1] = 24'b111111111010001110110001;
		character_jump[3][2] = 24'b000000000000000000000000;
		character_jump[3][3] = 24'b111111111010001110110001;
		character_jump[3][4] = 24'b000000000000000000000000;
		character_jump[3][5] = 24'b111111111010001110110001;
		character_jump[3][6] = 24'b000000000000000000000000;
		character_jump[3][7] = 24'b111111111010001110110001;
		character_jump[3][8] = 24'b000000000000000000000000;
		character_jump[3][9] = 24'b111111111010001110110001;
		character_jump[3][10] = 24'b111111111111001000000000;
		character_jump[4][0] = 24'b111111111010001110110001;
		character_jump[4][1] = 24'b111111111010001110110001;
		character_jump[4][2] = 24'b000000000000000000000000;
		character_jump[4][3] = 24'b111111111010001110110001;
		character_jump[4][4] = 24'b111111111010001110110001;
		character_jump[4][5] = 24'b111111111010001110110001;
		character_jump[4][6] = 24'b111111111010001110110001;
		character_jump[4][7] = 24'b111111111010001110110001;
		character_jump[4][8] = 24'b000000000000000000000000;
		character_jump[4][9] = 24'b111111111010001110110001;
		character_jump[4][10] = 24'b111111111010001110110001;
		character_jump[5][0] = 24'b111111111010001110110001;
		character_jump[5][1] = 24'b111111111010001110110001;
		character_jump[5][2] = 24'b000000000000000000000000;
		character_jump[5][3] = 24'b111111111010001110110001;
		character_jump[5][4] = 24'b111111111010001110110001;
		character_jump[5][5] = 24'b111111111010001110110001;
		character_jump[5][6] = 24'b111111111010001110110001;
		character_jump[5][7] = 24'b111111111010001110110001;
		character_jump[5][8] = 24'b000000000000000000000000;
		character_jump[5][9] = 24'b111111111010001110110001;
		character_jump[5][10] = 24'b111111111010001110110001;
		character_jump[6][0] = 24'b111111111010001110110001;
		character_jump[6][1] = 24'b111111111010001110110001;
		character_jump[6][2] = 24'b000000000000000000000000;
		character_jump[6][3] = 24'b000000000000000000000000;
		character_jump[6][4] = 24'b111111111010001110110001;
		character_jump[6][5] = 24'b111111111010001110110001;
		character_jump[6][6] = 24'b111111111010001110110001;
		character_jump[6][7] = 24'b000000000000000000000000;
		character_jump[6][8] = 24'b000000000000000000000000;
		character_jump[6][9] = 24'b111111111010001110110001;
		character_jump[6][10] = 24'b111111111010001110110001;
		character_jump[7][0] = 24'b111111111010001110110001;
		character_jump[7][1] = 24'b111111111010001110110001;
		character_jump[7][2] = 24'b111111111111111111111111;
		character_jump[7][3] = 24'b111111111010001110110001;
		character_jump[7][4] = 24'b111111111010001110110001;
		character_jump[7][5] = 24'b111111111010001110110001;
		character_jump[7][6] = 24'b111111111010001110110001;
		character_jump[7][7] = 24'b111111111010001110110001;
		character_jump[7][8] = 24'b111111111111111111111111;
		character_jump[7][9] = 24'b111111111010001110110001;
		character_jump[7][10] = 24'b111111111010001110110001;
		character_jump[8][0] = 24'b111111111010001110110001;
		character_jump[8][1] = 24'b111111111010001110110001;
		character_jump[8][2] = 24'b111111111111111111111111;
		character_jump[8][3] = 24'b111111111111111111111111;
		character_jump[8][4] = 24'b111111111010001110110001;
		character_jump[8][5] = 24'b111111111010001110110001;
		character_jump[8][6] = 24'b111111111010001110110001;
		character_jump[8][7] = 24'b111111111111111111111111;
		character_jump[8][8] = 24'b111111111111111111111111;
		character_jump[8][9] = 24'b111111111010001110110001;
		character_jump[8][10] = 24'b111111111010001110110001;
		character_jump[9][0] = 24'b000000000000000000000000;
		character_jump[9][1] = 24'b111111111010001110110001;
		character_jump[9][2] = 24'b111111111111111111111111;
		character_jump[9][3] = 24'b111111111111111111111111;
		character_jump[9][4] = 24'b111111111111111111111111;
		character_jump[9][5] = 24'b111111111010001110110001;
		character_jump[9][6] = 24'b111111111111111111111111;
		character_jump[9][7] = 24'b111111111111111111111111;
		character_jump[9][8] = 24'b111111111111111111111111;
		character_jump[9][9] = 24'b111111111010001110110001;
		character_jump[9][10] = 24'b000000000000000000000000;
		character_jump[10][0] = 24'b000000000000000000000000;
		character_jump[10][1] = 24'b000000000000000000000000;
		character_jump[10][2] = 24'b000000000000000000000000;
		character_jump[10][3] = 24'b111111111111111111111111;
		character_jump[10][4] = 24'b111111111111111111111111;
		character_jump[10][5] = 24'b111111111111111111111111;
		character_jump[10][6] = 24'b111111111111111111111111;
		character_jump[10][7] = 24'b111111111111111111111111;
		character_jump[10][8] = 24'b000000000000000000000000;
		character_jump[10][9] = 24'b000000000000000000000000;
		character_jump[10][10] = 24'b000000000000000000000000;
		character_jump[11][0] = 24'b000000000000000000000000;
		character_jump[11][1] = 24'b000000000000000000000000;
		character_jump[11][2] = 24'b000000000000000000000000;
		character_jump[11][3] = 24'b111111111111111111111111;
		character_jump[11][4] = 24'b111111111111111111111111;
		character_jump[11][5] = 24'b111111111111111111111111;
		character_jump[11][6] = 24'b111111111111111111111111;
		character_jump[11][7] = 24'b111111111111111111111111;
		character_jump[11][8] = 24'b000000000000000000000000;
		character_jump[11][9] = 24'b000000000000000000000000;
		character_jump[11][10] = 24'b000000000000000000000000;
		character_jump[12][0] = 24'b000000000000000000000000;
		character_jump[12][1] = 24'b000000000000000000000000;
		character_jump[12][2] = 24'b000000000000000000000000;
		character_jump[12][3] = 24'b111111111111111111111111;
		character_jump[12][4] = 24'b111111111111111111111111;
		character_jump[12][5] = 24'b111111111111111111111111;
		character_jump[12][6] = 24'b111111111111111111111111;
		character_jump[12][7] = 24'b111111111111111111111111;
		character_jump[12][8] = 24'b000000000000000000000000;
		character_jump[12][9] = 24'b000000000000000000000000;
		character_jump[12][10] = 24'b000000000000000000000000;
		character_jump[13][0] = 24'b000000000000000000000000;
		character_jump[13][1] = 24'b000000000000000000000000;
		character_jump[13][2] = 24'b000000000000000000000000;
		character_jump[13][3] = 24'b111111111111111111111111;
		character_jump[13][4] = 24'b111111111111111111111111;
		character_jump[13][5] = 24'b111111111111111111111111;
		character_jump[13][6] = 24'b111111111111111111111111;
		character_jump[13][7] = 24'b111111111111111111111111;
		character_jump[13][8] = 24'b000000000000000000000000;
		character_jump[13][9] = 24'b000000000000000000000000;
		character_jump[13][10] = 24'b000000000000000000000000;
		character_jump[14][0] = 24'b000000000000000000000000;
		character_jump[14][1] = 24'b000000000000000000000000;
		character_jump[14][2] = 24'b111111111111111111111111;
		character_jump[14][3] = 24'b111111111111111111111111;
		character_jump[14][4] = 24'b111111111111111111111111;
		character_jump[14][5] = 24'b111111111111111111111111;
		character_jump[14][6] = 24'b111111111111111111111111;
		character_jump[14][7] = 24'b111111111111111111111111;
		character_jump[14][8] = 24'b111111111111111111111111;
		character_jump[14][9] = 24'b000000000000000000000000;
		character_jump[14][10] = 24'b000000000000000000000000;
		character_jump[15][0] = 24'b000000000000000000000000;
		character_jump[15][1] = 24'b111111111111111111111111;
		character_jump[15][2] = 24'b111111111111111111111111;
		character_jump[15][3] = 24'b111111111111111111111111;
		character_jump[15][4] = 24'b000000000000000000000000;
		character_jump[15][5] = 24'b000000000000000000000000;
		character_jump[15][6] = 24'b000000000000000000000000;
		character_jump[15][7] = 24'b111111111111111111111111;
		character_jump[15][8] = 24'b111111111111111111111111;
		character_jump[15][9] = 24'b111111111111111111111111;
		character_jump[15][10] = 24'b000000000000000000000000;
		character_jump[16][0] = 24'b000000000000000000000000;
		character_jump[16][1] = 24'b111111111100000100000111;
		character_jump[16][2] = 24'b111111111100000100000111;
		character_jump[16][3] = 24'b111111111100000100000111;
		character_jump[16][4] = 24'b000000000000000000000000;
		character_jump[16][5] = 24'b000000000000000000000000;
		character_jump[16][6] = 24'b000000000000000000000000;
		character_jump[16][7] = 24'b111111111100000100000111;
		character_jump[16][8] = 24'b111111111100000100000111;
		character_jump[16][9] = 24'b111111111100000100000111;
		character_jump[16][10] = 24'b000000000000000000000000;
		character_jump[17][0] = 24'b000000000000000000000000;
		character_jump[17][1] = 24'b111111111100000100000111;
		character_jump[17][2] = 24'b111111111100000100000111;
		character_jump[17][3] = 24'b111111111100000100000111;
		character_jump[17][4] = 24'b000000000000000000000000;
		character_jump[17][5] = 24'b000000000000000000000000;
		character_jump[17][6] = 24'b000000000000000000000000;
		character_jump[17][7] = 24'b111111111100000100000111;
		character_jump[17][8] = 24'b111111111100000100000111;
		character_jump[17][9] = 24'b111111111100000100000111;
		character_jump[17][10] = 24'b000000000000000000000000;
	end
endmodule 